library verilog;
use verilog.vl_types.all;
entity Control_Unit_vlg_vec_tst is
end Control_Unit_vlg_vec_tst;
