library verilog;
use verilog.vl_types.all;
entity DEUARC_BUSYSTEM_vlg_vec_tst is
end DEUARC_BUSYSTEM_vlg_vec_tst;
